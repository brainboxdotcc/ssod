## Symtom:
Drabbade individer upplever en sjukt grön nyans på huden, åtföljd av ett gradvis förfall av kött. Trötthet, svaghet och allmän sjukdomskänsla är vanliga.

## Orsaker:
Dras samman genom exponering för vissa svampar som finns i fuktiga grottor och myrmarker. Sporer som frigörs av svamparna är det primära överföringssättet.

## Behandlingar:
En skicklig healer kan använda reningsbesvär för att rena kroppen från svampinfektionen. Sällsynta örter som finns i mystiska lundar kan användas i grötomslag för att underlätta återhämtningen.