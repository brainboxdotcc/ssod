Alver, höga och kungliga, står som majestätiska varelser utrustade med en djupgående behärskning av magi. Deras koppling till landet är helig, och betraktar det som en gudomlig gåva från gudarna. Alver vaktar våldsamt sina territorier, och varje försök att göra intrång på alvens domäner möts av snabbt fördömande, vilket stämplar inkräktarna som kättare.

Alvsamhället präglas av en djup respekt för auktoritet och ordning. Denna anslutning till hierarkin sträcker sig bortom militära sammanhang och sträcker sig in i själva familjelivet. I familjära miljöer intar fadern en ledarställning, och tomtarna följer plikttroget efter utan avvikande mening. Denna orubbliga lydnad är inte bara en fråga om tradition; det bottnar i en övertygelse om att faderns maktanvändning kommer att granskas i livet efter detta, ett heligt ansvar som inte får missbrukas.

Andlighet går genom alvernas ådror, och deras djupa förståelse för magi skiljer dem åt. De är medvetna om både dess välvilliga kapacitet och de potentiellt upprörande biverkningar den kan släppa lös. Magi blir en kanal för försvar, vilket gör det möjligt för dem att skydda sina hem, forma eteriska städer på himlen och till och med skymta en kort bit in i framtiden.

I Cryptillias intrikata gobeläng framträder alver som väktare av både det mystiska och det påtagliga. Deras engagemang för landets gudomliga helighet, deras disciplinerade hierarki och deras djupa koppling till den mystiska konsten bidrar till den gåtfulla och eteriska natur som definierar dessa lysande varelser och deras plats i världen.