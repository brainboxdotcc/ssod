Scythe Island, inbäddad i det tumultartade vattnet i Rushwatersundet, står som en ensam bastion i havet i de södra vidderna av Utopia. I hjärtat av denna mystiska ö ligger den förfallna Castle Scythe, en olycklig struktur höljd i rykten om ett mörkt och hemsökt förflutet. Slottet har varit övergivet i evigheter och utstrålar en luft av illvilja som gör det till ett oroande resmål för de modigaste äventyrare.

Själva omnämnandet av Castle Scythe framkallar berättelser om kusliga uppenbarelser, spöklika viskningar och oroande ekon från djupet av dess hemsökta salar. En gång i tiden ett säte för makt och auktoritet, står slottet nu som en spektral vaktpost som bevakar hemligheterna från en svunnen tid.

Legender talar om en härskare vars törst efter herravälde ledde till outsägliga illdåd inom slottets murar. Vissa hävdar att andarna hos de förorättade fortfarande dröjer kvar, utan att kunna finna vila. Andra viskar om eldgamla ritualer som utförs i slottets dolda kammare och lämnar efter sig en utomjordisk rest som genomsyrar luften.

Att närma sig Scythe Island möts av bävan, när den olycksbådande silhuetten av Castle Scythe skymtar vid horisonten. Många har vågat utforska dess ruiner och letat efter svar på de mysterier som omsluter det ödsliga slottet. Ändå är det få som återvänder med berättelser om sina fynd, och de som gör det talar i tysta toner om de oroande möten som väntar i Castle Scythes hemsökta salar. Ön står som ett skrämmande bevis på de kvardröjande skuggorna från dess förflutna, och lockar endast de djärvaste själarna att avslöja sanningen inom dess spektrala famn.