## Stava: Vatten

Med bara en gest frammanar vattenbesvärjelsen en strömmande ström från valfri del av kastarens form, som ofta gynnar handflatorna eller till och med ögonen för dramatisk känsla. Denna vattenkraft blir ett mångsidigt verktyg som tvingar fiender till ofördelaktiga positioner eller säkerställer överlevnad under svåra omständigheter, som att korsa en ödemark.