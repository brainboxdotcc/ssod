I den urbana gobelängen av Cryptillia, utspelar sig ett nät av fredsbevarande styrkor, känd som milisen, som en viktig tråd enligt kungligt dekret. Rikets herrar och damer är enligt lag bundna att samla dessa oberoende fredsbevarare, en styrka som är utformad för att upprätthålla ordningen i de livliga städerna och byarna. Det kungliga direktivet begränsar emellertid milisens uppgifter enbart till stadsområden, och anser att deras utplacering på landsbygden är en onödig utgift av tid och resurser.

Omfattningen och auktoriteten för varje milisenhet formas av den härskande herren eller damen i staden. Ändå framträder ofta en nyanserad verklighet under fredsbevarande fasaden. Många milisstyrkor, behäftade med korruption, befinner sig under kontroll av överordnade som prioriterar illusionen av att framgångsrikt bekämpa brottslighet framför äkta brottsbekämpning. Milisens motiv, som betalas per arresteringsbasis, kan luta mer mot ekonomisk vinning än strävan efter rättvisa. Förbered dig, för att möta lagens långa arm kan vara ett oundvikligt kapitel i din strävan, eftersom din arrestering kan fungera som en myntfylld välsignelse för männens plånböcker.

Beväpnad med tillstånd att utöva dödligt våld, arbetar milisen med ett omfattande mandat och tillämpar det inte bara på kända brottslingar utan även på misstänkta och de som gör motstånd mot arrestering. Konsekvenserna för överträdelser i Utopia och liknande länder är allvarliga, vilket främjar en miljö där brottsligheten begränsas och en bräcklig fred råder över städerna.

Ändå kan just den kraft som är avsedd att upprätthålla ordning ibland bli förebudet om oordning. Fall av milisuppror som lett till störtandet av rättmätiga herrar har registrerats. I sådana scenarier segrar ofta ändamålsenligheten, med kejsaren som förklarar den nye härskaren som den officiella herren, förutsatt att kungligt befallning upprätthålls. Den känsliga balansen mellan auktoritet och uppror formar berättelsen om milisen och målar upp en komplex bild av rättvisa, makt och strävan efter fred i Cryptillias urbana landskap.