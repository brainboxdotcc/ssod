I Cryptillias skuggiga underliv, ett rike där överlevnad ofta vacklar på gränsen till nödvändighet, finner en mängd invånare att de dras till ett liv i brott. Bland de olika nyanserna av överträdelse framträder tjuvar som de vanligaste, deras kvicka fingrar och hemliga färdigheter gör dem till kvintfigurerna i det kriminella landskapet.

Expertis i att få tillgång till säkrade domäner definierar tjuvarnas hantverk. Beväpnade med en intim förståelse för låsmekanismer navigerar dessa kvicka infiltratörer i tumblers intrikata dans med finessen hos erfarna hantverkare. Deras behärskning sträcker sig bortom det vardagliga och gräver ner i magins rike när de lär sig trollformler som "öppna", och reder ut hemligheterna som ligger bakom låsta dörrar.

Stealth blir en andra natur för tjuvar, deras rörelser höljda i tystnadens och bedrägeriernas slöjor. Bortom låsplockningens rike har många finslipat sina färdigheter i den hemliga konsten att plocka i fickorna, navigera på trånga gator med en nästan kuslig förmåga att befria värdesaker utan att väcka misstankar.

Tjuvar är dock inte begränsade till skuggorna enbart för skändliga syften. Deras smidighet och list gör dem till exceptionella scouter, kapabla att glida förbi hårt bevakade utposter med fantomernas finess. I stridens kaos förvandlar deras förmåga att infiltrera, samla intelligens och slå snabbt från oväntade vinklar dem till värdefulla tillgångar.

Under faner av uppenbar knapphet samlar tjuvar ofta stora rikedomar. Deras list och påhittighet tillåter dem att avslöja dolda skatter, vilket vänder oddsen till deras fördel. Alltså, vad som kan tyckas vara en ödmjuk tillvaro döljer den subtila överflöden hos dem som är skickliga på att manövrera genom den invecklade väven i Cryptillias kriminella landskap.