Demoner manifesterar sig inom Cryptillia som ett påtagligt och bevisat hot, existerande som enheter av ren energi med den unika förmågan att materialisera sig efter behag. Dessa uråldriga varelser är före ankomsten av människor och orcher, som går tillbaka över tre årtusenden, och deras eteriska rike är naturligt knutet till ursprunget till magi och förekomsten av magiska artefakter i Cryptillia.

Demoner hyser ett djupt förakt och hat mot varelser som är bundna av fysisk materia och anser dem vara underlägsna. Deras intelligens, som vida överträffar dödliga varelsers, har lett dem att korsa inte bara Cryptillias vidd utan även de omgivande stjärnsystemen, utan hinder av ömtåliga miljöer som begränsar människor.

För att utöva ett betydande inflytande på den fysiska världen, genomför demoner en komplex process. De måste äga en fysisk varelse genom att kartlägga sin energi i samma neurala mönster som en humanoid varelse, vilket effektivt skriver över det befintliga medvetandet. Denna komplicerade procedur kräver tid, ansträngning och precision, vilket ofta kräver en distraktion, som en ceremoni eller en långvarig trollformel. Synkroniseringen med värdens kropp, avgörande för att upprätthålla viktiga funktioner som hjärtslag, gör sömnen till ett lämpligt ögonblick för denna kosmiska invasion.

När den lyckas tar demonen kontroll över värdens fysiska kropp och utrotar alla spår av den förra varelsen. Den manipulerade varelsen blir sedan ett instrument för att skapa förödelse i den fysiska världen, och rensa vägen för demoner att återta Cryptillia som de hade gjort i miljontals år innan mänsklighetens ankomst.

Endast de mäktigaste trollkarlarna förstår allvaret i detta existentiella hot mot allt fysiskt liv. Deras medvetenhet får dem att utfärda varningar till dem som har tillräckligt med intelligens för att förstå faran, och samlar i hemlighet en hemlig armé som förberedelse för den oundvikliga dagen då domen faller över Cryptillia. Det hotande hotet om demonisk besittning, dolt i skuggorna, understryker den känsliga balansen mellan den magiska och fysiska världen i denna fantastiska värld.