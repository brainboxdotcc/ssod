Hartleaf, en delikat ört som frodas i de bördiga jordarna i Cryptillia, är sammanflätad med essensen av rörelse och vatten. Dess smala stjälkar, prydda med hjärtformade löv, skimrar med ett subtilt akvatiskt sken. När den skördas under silverljuset från en halvmåne, sägs örtens styrka nå sin zenit. Trollkarlar och trollkastare prisar Hartleaf för dess koppling till smidighet och snabbhet, och använder den ofta som en nyckelkomponent i trollformler som åberopar smidiga rörelser eller manipulerar vattenströmmar.