The First Age of Magic är en period av tidig kryptillian historia som framstår som en skugg epok, en era höljd i tidens dimmor när hela världen var snärjd i en utdragen magisk konflikt som varade i århundraden. Det var en period som föregick upplysningen av många raser om trollformningens farliga natur, en tid då den verkliga omfattningen av det demoniska hotet, som lurar i de osynliga energierna kring Cryptillia, förblev beslöjade.

Konflikten varade tills ett avgörande ögonblick då flera visionära trollkarlar slöt en aldrig tidigare skådad allians, överskridande gränserna som en gång hade ställt alver, människor och dvärgar mot varandra. Förenade i syfte orkestrerade de ett historiskt fredsavtal, en pakt etsad med magins kraftfulla trådar i ett försök att väva en bestående fred i århundraden, om inte evigheten.

Det eteriska bläcket på detta magiska pergament var dock inte torrt innan dess brister visade sig. Ilska krafter, som tros vara demoners intrig, ingrep med skändlig avsikt, omintetgjorde rasernas enhet och hindrade vissa från att delta i fredstoppmötet. Särskilt frånvarande var Orc-imperiet och vissa alverstammar, ödesbestämda att avvika in i den olycksbådande härstamningen som kallas mörkalverna.

Frånvaron av dessa raser från fredspakten introducerade en irreparabel spricka i strukturen av den föreställda eviga freden. Den olycksbådande agendan som dessa utestängda raser hade, försökte inte bara utplåna de ideal som inkapslades i fredspakten utan också att avveckla själva upprätthållarna av fördraget. Spöket av ständiga konflikter dröjde sig kvar och kastade en lång skugga över de utopiska strävanden i ett rike som längtade efter en bestående fred som för alltid verkade svårfångad.

I den kryptilliska historiens gobeläng står Magins första tidsålder som en varnande berättelse, en krönika som ekar med konsekvenserna av okontrollerad magisk kraft, demoniskt inflytandes bedrägeri och pakternas bräckliga natur som är avsedda att binda en splittrad värld.