Wizards Ivy, en växt höljd i mystik och vördad för sina djupa magiska egenskaper, trivs i de dolda hörnen av Cryptillia. Sällsynt och svårfångad, sägs denna murgröna ha oöverträffad magisk energi. Trollkarlar och arkanister eftertraktar det för dess potential att förstärka spellcasting-förmågor. När de är noggrant integrerade i trollformler, fungerar Wizards Ivy som en katalysator och förstärker de mystiska energierna som kanaliseras av kastaren. Växtens invecklade vinstockar och självlysande löv antyder en koppling till uråldriga mystiska krafter, vilket gör den till en eftertraktad komponent i jakten på magiskt mästerskap.