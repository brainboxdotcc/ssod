## Stava: Vapenfärdighet

Vapenfärdighetsbesvärjelsen, som liknar den svårfångade dansen av "smyga" besvärjelsen, påverkar trollkarlens stridsfinesser. Vid anropet genomgår kastarens skicklighetspoäng en spektakulär fyrdubbling, vilket gör dem till en formidabel kraft på slagfältet under en varaktighet av fem stycken. Efterdyningarna är dock en övergående svacka, eftersom skicklighetspoängen sjunker till hälften av sitt ursprungliga värde under en motsvarande varaktighet. Dessa effekter ackumuleras med successiva spellcasting, vilket kräver ett strategiskt tillvägagångssätt för att frigöra den fulla potentialen hos denna stridscentrerade förtrollning.