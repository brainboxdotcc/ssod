Port Obligan, inbäddat längs Utopias södra stränder, står som en livlig hamnstad och en viktig inkörsport till Rushwatersundet. Detta strategiska läge gör det till ett viktigt handelsnav för de södra regionerna på kontinenten, vilket underlättar utbyte av varor, kunskap och kultur.

När fartyg kommer och går skapar de rytmiska ljuden av vågor och avlägsna måsar en symfoni längs de livliga hamnen. Hamnen är livlig med aktivitet, med en blandning av lastfartyg, handelsfartyg och örlogsfartyg som navigerar i Rushwatersundet.

Arkitekturen i Port Obligan är en blandning av funktionalitet och maritim charm. Stabila lager kantar vattnet och lagrar varor på väg till avlägsna länder. Tavernor och värdshus vänder sig till sjömän och handlare och erbjuder andrum och kamratskap. Den salta brisen bär doften av havet och blandas med handelns livliga energi.

Stadens gator är en labyrint av kullerstensvägar som leder till olika marknadsplatser, skråhallar och bostadskvarter. Köpmän säljer sina varor på livliga marknader, medan hantverkare finslipar sina kunskaper i verkstäder utspridda över hela staden.

Trots dess ekonomiska betydelse står Port Obligan inför ett ständigt närvarande hot från den närliggande Demon Lord Garneths befästa borg. Den olycksbådande silhuetten av Garneths fäste skymtar i fjärran, en ständig påminnelse om den osäkra balansen mellan handel och det lurande mörkret.

Staden har en påtaglig luft av motståndskraft, eftersom dess invånare förstår den känsliga dansen mellan välstånd och fara. Den lokala milisen håller ett vakande öga på horisonten, redo att försvara sig mot alla inträngande hot. Trots det hotande hotet fortsätter Port Obligan att frodas som ett avgörande maritimt centrum, som navigerar i det ömtåliga vattnet mellan handeln och skuggan av Garneths fäste.