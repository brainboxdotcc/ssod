Elfbane, en eterisk ört som blomstrar i närheten av snabbrörliga fåglar, väver sina rötter djupt i luftens mystiska energier. Örtens smala grenar bär känsliga, fjäderliknande löv som prasslar med ekon av fågelvindar. Legender talar om Elfbanes förtrollande lockelse och hämtar inspiration från fåglarnas snabbhet i flykt. Spellcasters skickliga i kryptillianflorans krångligheter införlivar ofta Elfbane i sina hopkok, och tror att dess essens förstärker trollformler relaterade till snabbhet, grace och de luftiga rikena.