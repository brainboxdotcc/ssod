## Stava: Styrka

Styrkebesvärjelsen, en flyktig våg av onaturlig styrka, ger kastaren omänsklig styrka under en bråkdel av tiden. Vanligtvis utnyttjas i de kortaste intervallen, det ger kastaren möjligheten att släppa lös ett förödande slag mot en motståndare, vilket får dem att slingra sig från den överväldigande kraften.