## Stava: Sköld

Shield-besvärjelsen, en bastion av magiskt försvar, frammanar en skyddande bubbla som omsluter kastaren och potentiella allierade. Denna eteriska barriär har en rustningspoäng på 6 och håller i tio spelstycken. Dess tillämpning är dock beroende av tillgången till en betydande period av ledig tid för casting. Att försöka åberopa denna besvärjelse i striden, med motståndare som närmar sig, är oklokt. En försiktig kastare reserverar sin användning för stunder av strategiska fördelar under perioder av andrum.