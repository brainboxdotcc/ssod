Guldslätten, som sträcker sig så långt ögat kan se i de södra delarna av Cryptillia, presenterar en spökande och ödslig tablå. En gång i tiden ett landskap som kan ha blomstrat med mångsidigt liv, bär regionen nu ärren av en gammal katastrofal händelse. Det verkar som om själva landet har "glasat", som om någon illvillig kraft hade skrivit över den naturliga ordningen.

I denna vidsträckta vidd av ödslighet, där livet kämpar för att slå rot, står Port Krellis magra tillvaro. Den här kuststaden ligger inbäddat längst ut i södra delen av landet och håller fast vid överlevnaden genom att utnyttja havets rikedom. Dess motståndskraftiga invånare, beroende av havets överflöd, har anpassat sig till sina tuffa omgivningar och fått ett blygsamt liv mitt i de oförlåtande guldslätterna.

Nära Port Krellis ligger en dyster påminnelse om regionens farliga natur - Nattugglans vrak. Fartyget var en gång en majestätisk galjon och dukade under för de häftiga elementen under en kraftig storm för många år sedan. Nu ligger skelettresterna av fartyget utspridda längs kusten och fungerar som både en gripande symbol för det oförutsägbara havet och ett bevis på de utmaningar som de som trotsar Cryptillias vatten står inför. Resterna av Nattugglan står som ett tyst vittne till de formidabla krafter som formar ödet för detta ödsliga och krossade land.