## Symtom:
Svullna, smärtsamma lymfkörtlar (buboer), hög feber, frossa och trötthet. I svåra fall leder det till septikemi och organsvikt.

## Orsaker:
smittats av infekterade loppor, som ofta angriper gnagare. Vanlig i trånga stadsområden och regioner med dålig sanitet.

## Behandlingar:
Reningsbesvär kan hjälpa till att bekämpa infektionen. Den sällsynta Starpetal-örten, som finns i avlägsna bergsregioner, tros ha potenta antibakteriella egenskaper.