## Symtom:
Snabb försämring av blodkärlen, vilket orsakar inre blödningar, svår anemi och organsvikt. Mörkt, nästan svart blod är en distinkt egenskap.

## Orsaker:
Smittas genom bett av infekterade varelser eller genom kontakt med kontaminerat blod. Vanligt i områden där mörk magi är utbredd.

## Behandlingar:
Magiska helande besvärjelser fokuserade på blodrening kan bromsa utvecklingen. Extrakt från Silvermoon-blomman, som finns i heliga trädgårdar, har känt till att motverka effekterna.