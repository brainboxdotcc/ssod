Hallucinogen, en kraftfull ört som frodas i de vilda och otämjda hörnen av Cryptillia, har kraften att förändra uppfattningar för dem som tar del av dess väsen. Hallucinogen känns igen på sina livfulla, mångfärgade blommor och är eftertraktad av shamaner och illusionister för sina hallucinatoriska egenskaper. När det integreras i trollformler framkallar Hallucinogen en tillfällig avvikelse från verkligheten, vilket gör att de inom dess inflytande upplever levande och förvrängda syner. Den utövas av trollformler som försöker desorientera motståndare eller utforska förändrade medvetandetillstånd.