## Stava: E.S.P.

E.S.P., en kanal till sinnets fördjupningar, tillåter en kastare att fördjupa sig i tankar, implantera illusioner som styr fiender mot självförvållad skada eller oavsiktliga fördelar. Dess styrka, besläktad med hypnotism, finner sin värld utanför stridens kaos. Genom att utnyttja sårbarheterna hos ett ofokuserat och svagt sinne, E.S.P. uppenbarar strategiska fördelar i subtilare engagemang, strategiska manipulationer och den subtila dansen av intelligens. I händerna på en klok trollkarl, E.S.P. avslöjar den intrikata väven av avsikter, förvandlar slagfältet till ett skede av mentalt schack.