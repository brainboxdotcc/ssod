I de avlägsna ekona av kryptillians historia samlades en koalition av raser för att upprätta den legendariska "fredspakten". Ledare från olika världar, inklusive det mänskliga imperiet, alfstammarna och dvärgarna, samlades med den ädla avsikten att inviga en era av harmoni över hela planeten. Emellertid, mitt i denna monumentala församlings storhet, insinuerade sig en skändlig korruption, som kastade en skugga över strävan efter enhet.

När de stora fredsfartygen seglade över Stora havets vidd, på väg mot de neutrala länder som valts ut för det avgörande mötet och undertecknandet av pakten, ingrep mörka krafter. Osynliga och illvilliga avbröt dessa krafter den fridfulla resan och avledde flera fartyg ur kurs med stormar, konstiga monster och andra onaturliga fenomen. Tyvärr, den avsedda destinationen vid stranden av den utsedda ön bevittnade frånvaron av många armadas, för alltid förlorade till de oförutsägbara nyckerna från den mystiska störningen.

Bland de olyckliga offren för detta förvrängda öde fanns en hel alvstam, avskild från de magiska skydd som utlovades av fredspakten. Isolerade och övergivna hyste alverna förbittring, en känsla som växte fram med tiden. Utan paktens mystiska sköld växte de till att förakta de ideal den symboliserade, och vände sig slutligen mot själva magin som försökte bevara den bräckliga freden i Cryptillia. Denna en gång ädla alvstam förvandlades till "Mörka alverna".

De mörka alverna, nu befläckade av misstro och fiendskap mot utomstående, övergav principerna för öppen förhandling. De föredrog skuggor framför ljuset och antog ett listigt tillvägagångssätt och lurade i bakgrunden för att observera världen obemärkt. Deras affärer blev präglade av bedrägeri, och de mörka underströmmar som de introducerade undergrävde magin som var avsedd att skydda rikets osäkra lugn.

Idag representerar mörkalverna opålitlighet och hat, deras handlingar är ett konstant hot mot den känsliga balansen som upprätthålls av resterna av fredspakten. Med en förkärlek för tyst manipulation och en preferens för förräderi framför öppen diskurs, navigerar Dark Elves i Cryptillias invecklade nät av allianser och fientligheter, och lämnar ett outplånligt märke på den ständigt utvecklande gobelängen i denna fantastiska värld.