I de olika länderna i Cryptillia har flera religioner utvecklats som en återspegling av deras tumultartade upplevelser och interaktioner med de magiska krafter som formar deras värld. De rådande trossystemen formas av historiska händelser, möten med mystiska enheter och den pågående kampen mellan ljus och mörker.

## The Church of the Arcane Light
Church of the Arcane Light, som grundades i efterdyningarna av den första tiden av magi, vördar de välvilliga aspekterna av magi. Anhängare tror på en gudomlig kraft som förkroppsligar den harmoniska balansen av magiska energier. De ser magi som en gåva från högre världar, skänkt till dödliga för att åstadkomma välstånd och upplysning. Prästerskapet, känt som Illuminators, strävar efter att utnyttja magiska energier för att förbättra samhället och för att bekämpa mörkrets krafter.

## Orden för evig vaksamhet
Född ur de obevekliga konflikterna med demoniska enheter, är Order of Eternal Vigilance en krigsreligiös orden. Dess anhängare, kända som Sentinels, ägnar sig åt att skydda mänskligheten från demoniska intrång. De tror att kampen mot mörka krafter är en evig strävan och att det krävs evig vaksamhet för att skydda rikena. Ritualistiska ceremonier involverar rening av vapen och skandering av uråldriga besvärjelser för att stärka barriärerna mellan världar.

## Sökarna av den dolda vägen
En mystisk och esoterisk sekt, Sökarna av den dolda vägen gräver ner sig i mysterierna med forntida rullar och bortglömda kunskaper. De vördar de magiska artefakterna som är utspridda över Cryptillia, och anser att de är nyckeln till att låsa upp djupare sanningar. De trogna, kallade sändebud, ger sig ut på uppdrag för att avslöja dold kunskap och dechiffrera de gåtfulla profetiorna som formar deras öde. Sökarna tror att upplysning ligger i att förstå de mystiska mysterier som vävts in i verklighetens väv.

## The Wayfarers' Fellowship
För dem som omfamnar den nomadiska livsstilen och navigerar i farorna med Cryptillias olika landskap, erbjuder Wayfarers' Fellowship tröst. Tillägnad resenärernas skyddsgud, betonar denna religion anpassningsförmåga och fyndighet. Pilgrimsfärder involverar att korsa förrädiska terränger och hylla heliga landmärken som tros innehålla gudomens väsen. Wayfarers tror att deras gudom vägleder dem genom livets ständigt föränderliga vägar.