Spikegrass, en motståndskraftig och farlig växt utspridda i Cryptillias farliga landskap, har knivskarpa blad som gör den till en formidabel trollformningskomponent. Växtens särdrag är dess sågtandade blad som liknar finslipade blad. Spellcasters med en förkärlek för offensiva förtrollningar gynnar Spikegrass, och använder dess naturliga skärpa för att förstärka trollformler som är utformade för att skära igenom magiska barriärer eller orsaka exakt skada. När det ingjuts i besvärjelser, ger Spikegrass sin spets till de mystiska krafterna som spelar, vilket förstärker besvärjelsens styrka och precision.