I det mystiska riket Cryptillia ger sig trollkarlar ut på en mödosam resa och ägnar större delen av sina liv åt att nysta upp den invecklade väven av magiska trollformler och trolldrycker. Magi här är inte ett privilegium reserverat för de få utvalda; snarare är det en latent förmåga som är inneboende i varje varelse. Men att behärska dessa magiska gåvor kräver år av orubblig övning, meditation och en djupgående förståelse för farorna som lurar inom spellcasting.

Magi, i sin essens, hämtas från de omgivande energierna som omsluter omgivningen. Processen med spellcasting involverar skicklig manipulation av rå energi – oavsett om det är värmen som kommer från en flammande eld eller den kinetiska energin som härrör från rörelse. Trollkarlens sinne fungerar som kanalen och formar dessa energier till en mer målmedveten och kontrollerad form. Förvecklingarna i denna transformativa process förblir höljda i mystik, en gåta som fängslar de nyfikna sinnena hos Cryptillias invånare.

Mitt i detta magiska landskap trotsar vissa varelser tillvarons konventionella regler. Demoner och eteriska uppenbarelser, till exempel, verkar på en metabolism som drivs helt av energi. Dessa entiteter, drivna av sin illvilliga natur, har förmågan att överföra sina energier till materiebaserade varelser. Konsekvensen är besittning, en farlig handling som ger demonen fullständig kontroll över värden. I fallet med en guide kan detta intrång visa sig vara mycket farligt, vilket ofta resulterar i förödande resultat.

När trollkarlar beträder den känsliga balansen mellan att utnyttja energierna runt dem och att skydda sig själva från de rovdjur som dras till deras makt, blir den mystiska konsten både en källa till vördnad och bävan i Cryptillia. I jakten på magiskt behärskning navigerar trollkarlar i det okända och gräver ner sig i mysterierna som ligger till grund för själva strukturen i deras mystiska tillvaro.