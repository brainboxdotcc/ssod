## Förtrollning: Woodsmanship

Woodsmanship-förtrollningen, en harmonisk blandning av naturens väsen och mystiska behärskning, förlänar för ett ögonblick kastaren med en skogsmans omfattande färdigheter. Denna förtrollande infusion sträcker sig inte bara till den invecklade kunskapen om skogsmarker utan integreras sömlöst med gjutmaskinens befintliga skicklighet. Besvärjelsens inflytande sträcker sig över exakt en dag och erbjuder en övergående men ändå uppslukande koppling till den sylviska konsten. Men att anpassa sig till sådan skogsskicklighet kräver en tålmodig cykel, vilket tillåter att besvärjelsen bara kan kastas en gång varje spelvecka.