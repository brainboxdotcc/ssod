I Cryptillias tumultartade sfärer dyker orker fram som en obeveklig kraft, som förkroppsligar en grymhet som återkommer genom varje handling. Våld är deras folkspråk, förhandling ett främmande begrepp eftersom de gynnar stridens trubbiga kraft framför dialogens nyanser. Med ett språk som ekar i gutturala toner och en upplevd lägre nivå av intelligens, organiserar orker sig i stamstrukturer, var och en styrd av en krigsherre flankerad av en kader av rådgivare, handplockade av krigsherren själv.

Även om det är teoretiskt accepterat att krigsherren bör lyssna till dessa rådgivares råd, beror verkligheten ofta på krigsherrens nyckfulla nycker. Orcher, drivna av sin inneboende stridbara natur, tillbringar större delen av sin existens i stridens strid. I avsaknad av en lämplig extern motståndare vänder de sig mot sig själva i en obeveklig cykel av inbördes konflikter. Vapenkollisionen och aggressionens dån definierar rytmen i deras dagliga liv.

När de inte är nedsänkta i strid, övergår orker mellan perioder av vila och fest, och njuter av efterdyningarna av sina erövringar. Galt- eller hästkött är basen i deras köttätande festmåltider, kompletterat med allt annat kött som kommer inom deras räckhåll. Den orchiska livsstilen blir en oändlig cykel av brutalitet, som växlar mellan stridens kaos, återställande slumrande och frossande fest.

Ett visceralt förakt definierar den orchiska uppfattningen av alver, en fiendskap som bottnar i ett djupt hat mot den naturliga världens alvervördnad. Om de fick valet att släppa lös sin aggression mot vilken ras som helst, skulle orker utan tvekan rikta in sig på alver, intensiteten av deras fiendskap påtaglig. Dvärgar, deras näst mest avskyvärda motståndare, delar en djupt rotad fiendskap som går tillbaka till magins tidigaste åldrar. I ett fruktansvärt kapitel av historien fördrev forntida dvärgar med tvång de ursprungliga orchiska invånarna från deras förfäders hemland, vilket antände en fejd som har bestått genom tiderna.

I Cryptillias vilda landskap står orcher som ett formidabelt bevis på aggressionens ohämmade kraft och ett hat som sträcker sig över generationer. Deras krigiska natur, stamsamhällen och bloddränkta historia sätter ett outplånligt märke på tapeten av den fantastiska värld de lever i.