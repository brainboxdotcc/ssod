## Stava: Ljus

En strålande aura materialiserar sig ovanför kastarens huvud med den lätta besvärjelsen, som ger en briljans som konkurrerar med alla lyktor. Denna förtrollade belysning trotsar att släcka om inte kastaren ger efter för att besegra eller avsiktligt drar tillbaka besvärjelsen, vilket ger en konstant källa av strålande utstrålning i de mörkaste världarna.