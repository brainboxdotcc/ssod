## Stava: Väx

Grow-förtrollningen, en motpol till dess krympande motsvarighet, åberopar utvidgningen av castern till proportioner begränsade endast av deras mystiska skicklighet. Denna formförstoring tjänar som en strategisk fördel, och ger trollkarlen större fysisk närvaro och, till synes, ökad skicklighet. Den försiktige utövaren måste dock utöva urskillning när han väljer det lämpliga ögonblicket för besvärjelsens avslutning, speciellt när den är omringad av höga fiender. Den mystiska förstärkningen, även om den är formidabel, kräver omdömesgill övervägande för att undvika oavsiktliga konsekvenser och säkerställa att kastaren sömlöst återintegrerar i den naturliga ordningen i sin miljö.