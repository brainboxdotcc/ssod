# Symtom:
Ihållande hosta, andningssvårigheter och ett raspande ljud vid inandning. Drabbade individer lider av försvagad lungfunktion och kan utveckla lunginflammation.

## Orsaker:
Inandning av luftburna sporer som frigörs av vissa giftiga växter och svampar som finns i mörka skogar. Exponering beror ofta på långvarig vistelse i sådana miljöer.

## Behandlingar:
Läkande besvärjelser som stärker andningsfunktionerna kan hjälpa till att återhämta sig. Den sällsynta Moonshade-örten, odlad i specifika alkemiska trädgårdar, är känd för sin kraft vid behandling av lungrelaterade sjukdomar.