I det vidsträckta riket Utopia står den ökända Demon Garneth som den mest formidabla motståndaren, en skugga som skymtar inte bara över den södra vidden utan kastar en mörk slöja över hela Cryptillia. En gång en mäktig herre som höll herraväldet över en stor del av södra Utopia, blev Garneths nedgång till illvilja ett spökande kapitel i landets historia.

I tidens annaler berättas det att Lord Garneth, driven av en omättlig makttörst och en begärlig önskan att utöka sitt territoriella domän, gav efter för ondskans lömska krafter. Den exakta katalysatorn för hans korruption förblir höljd i mystik, förlorad till tidernas viskningar. Hans en gång så storslagna slott, som nu var ett olyckligt fäste, blev en bastion av mörker, vars murar dolde den illvilliga herre som barrikaderade sig inombords.

Under ett halvt sekel har Garneths demoniska inflytande vuxit, spridit sig som ett elakartat nät och fångat landet i rädsla. Ingen levande själ har sett Lord Garneth sedan tiden för hans innehav, hans fysiska närvaro begränsad till slottets förbannade djup. Den en gång så välmående regionen under hans styre har blivit en förbjuden zon, en plats där ingen vågar beträda.

Även om Garneth själv förblir svårfångad, strövar hans hantlangare, förkroppsliganden av terror, fritt och sprider sin illvilja över landet. Från Larret-bron i norr till den livliga hamnstaden Port Obligan i söder, sträcker sig rankorna av hans inflytande långt och brett och lämnar ett spår av förtvivlan i deras spår.

Genom åren har berättelsen om Garneths skräckvälde etsat sig fast i Utopias kollektiva medvetande. Ändå, trots de otaliga skräckhistorierna och den utbredda kunskapen om hans illvilja, har ingen kommit fram med modet att konfrontera Garneth och få ett slut på hans tyranniska styre. De olycksbådande skuggorna av slottet står fortfarande kvar, och utmaningen att möta Garneth i en sista konfrontation väntar på en hjälte som är modig nog att kliva fram i den episka kampen mot mörkret som omsluter riket.