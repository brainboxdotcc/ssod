Stickwart, en sällsynt ört med gåtfulla ursprung, är genomsyrad av berättelser om telepatisk skicklighet. Inbäddat i de avlägsna delarna av Cryptillia, tros denna ört ha den extraordinära förmågan att ge användarna insikter i andras tankar. Trollkarlar och tankefokuserade spellcasters söker ofta efter Stickwart för dess påstådda tankeläsande egenskaper. När den ingår i trollformler, fungerar Stickwart som en kanal, förhöjer kastarens mentala skärpa och underlättar en kort gemenskap med de innersta tankarna hos dem i närheten.