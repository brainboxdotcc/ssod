## Stava: Eld

Eldbesvärjelsen, en dans av kontrollerade lågor på kastarens fingertoppar, förvandlar erfarna användare till utövare av eldstyrka. Mästare kan släppa lös det som en eldkastare, förvandla elementet till ett skräckinjagande vapen mot motståndare eller en tröstande källa till värme, en ledstjärna i kylan.