I historiens enorma annaler framträder barbarer som en uråldrig avvikelse från mänskligheten, och utvecklas under årtusenden av isolering till ett distinkt samhälle med sina egna övertygelser, teknologier och seder. Det är först under de senaste åren som dvärgforskare har avslöjat den avskilda existensen av barbarisk art i de kyliga delarna av de långt norra ödena i Cryptillia.

Mötet med dvärgarna var ett avgörande ögonblick för barbarerna, eftersom de flitiga upptäcktsresandena tillhandahöll ovärderlig kunskap och verktyg för att navigera i den hårda nordliga miljön. I kölvattnet av denna upptäckt har en våg av barbariska upptäcktsresande vågat sig söderut, ivriga att på egen hand bevittna de underverk och fristaden som kännetecknar det stora mänskliga imperiet.

På grund av sin långvariga isolering befinner sig barbarer avlastade av komplexa allianser och fiendskap. I allmänhet förkroppsligar de neutralitet, förtroende och en mottaglig natur, vilket gör dem lätta att delta i förhandlingar. Den enorma tid som spenderats i avskildhet har främjat en genuin nyfikenhet och öppenhet bland barbarerna, när de navigerar i komplexiteten i de "nya" länderna söderut, och söker förståelse och koppling till den expansiva mänskliga civilisationen.

När gränserna mellan kulturer suddas ut och ekon av uråldrig isolering bleknar, står barbarerna vid tröskeln till en ny era, redo att knyta förbindelser och bygga allianser med de olika samhällena som befolkar Cryptillia. Neutraliteten som definierar dem blir en bro, en grund på vilken nya relationer kan konstrueras, och den outnyttjade potentialen hos barbariska arter vecklas ut i den utspelade gobelängen av den mångfaldiga och dynamiska värld de nu utforskar.