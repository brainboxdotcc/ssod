Eldfrön, en kraftfull ört som frodas i de tempererade områdena i Cryptillia, är naturligt knuten till de ursprungliga krafterna av värme och eld. Denna anmärkningsvärda ört bär brinnande röda blommor som liknar miniatyrlågor och utstrålar värme även i de kyligaste miljöer. Trollkarlar och pyromaner omhuldar Fireseeds som en avgörande komponent i trollformler som utnyttjar de brinnande energierna i det mystiska. Fröna, när de krossas eller antänds under gjutningsprocessen, släpper lös en våg av intensiv värme, vilket förstärker glöden hos brandbaserade besvärjelser.