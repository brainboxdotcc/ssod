Blidvines, en mystisk ört gömd i de skuggiga hörnen av Cryptillia, är vördad för sin förmåga att avslöja dolda sanningar och dolda verkligheter. Vinrankorna, prydda med eteriska, självlysande blommor, verkar pulsera med ett utomjordiskt sken. Spellcasters som försöker reda ut mysterier eller avslöja de osynliga gynnar Blidvines som en viktig ingrediens i deras magiska brygger. När Blidvines ingjuts i besvärjelser, fungerar Blidvines som en metafysisk lykta, som lyser upp det mörka och avslöjar hemligheterna gömda i verklighetens veck.