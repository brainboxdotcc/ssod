## Valley City regional karta