Woodweed, en mångsidig ört som finns i hjärtat av Cryptillia, har unika egenskaper som underlättar snabba förändringar i storlek. Dess trådiga stjälkar och fjädrande blad anpassar sig sömlöst till fluktuationer i magiska energier. Trollkarlar som försöker manipulera dimensioner och ändra fysiska proportioner vänder sig ofta till Woodweed som en avgörande trollkastningskomponent. När den är noggrant integrerad i besvärjelser, gör Woodweed det möjligt för kastaren att korsa storleksmanipulationens världar med finess, vilket ger dem behärskning över ebb och flöde av rumsliga dimensioner.