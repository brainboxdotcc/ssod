Stava: Bolt

En manifestation av destruktiv styrka, bultförtrollningen driver fram en brännande, överhettad plasmabult från hjulets fingertoppar. Även om den är distinkt i sina effekter, förtjänar denna mystiska urladdning sin moniker som "lillebror" till trollformelns besvärjelse, med formidabel kraft och formidabla detaljer som utmärker den i riket av magiska projektiler.