Goblins är en motståndskraftig men ändå förslavad ras, fjättrad av orkstammarnas herravälde. Karaktäriserad av begränsad intelligens, troll har en kvick läggning som gör dem skickliga på att utföra enkla uppgifter, vilket gör dem till det föredragna valet framför mindre orcher för snåla uppgifter som att ta hand om galtar och skicka tillfångatagna hästar för de hemska stridsbanketter som markerar deras existens.

Goblins hyser ett kalkylerande men rättframt tänkesätt. Deras uppfinningsrikedom blir, när de slås samman, en gnista som kan antända uppror. När flera troll samarbetar överskrider deras kollektiva påhittighet deras individuella begränsningar, vilket gör det möjligt för dem att störta sina Orc-övervakare i massor. I en vågad revolt kan de svärma ut ur fångenskapens gränser och söka frihet och ett eget liv mitt i den otämjda vildmarken.

Trots sin ringa storlek, motsvarande den hos dvärgar, använder troll ett begränsat utbud av vapen. Men deras storlek motsäger deras motståndskraft i strid. Gäckande och smidiga, troll visar sig vara anmärkningsvärt utmanande mål som undviker sina motståndares strejker med otrolig skicklighet. I stridens närstrid blir deras kvickhet ett kraftfullt försvar, som kompenserar för deras blygsamma vapen med en undvikande skicklighet som frustrerar dem som försöker betvinga dem.

När troll navigerar i den förrädiska terrängen av träldom, uppror och den otämjda vildmarken, representerar de den okuvliga ande som kvarstår inför förtrycket. Deras berättelser väver en berättelse om listig överlevnad, samarbetsuppror och en motståndskraft som motsäger deras förslavade status i Cryptillias fantastiska gobeläng.