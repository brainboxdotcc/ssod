## Stava: Stjäla

Stjälbesvärjelsen, en flyktig åberopande av stöld, ger kastaren möjlighet att dubbla sin smygpoäng under en kort period. Besvärjelsens effekter kvarstår under ett enda spelstycke, följt av en obligatorisk nedkylning av tio stycken på grund av dess invecklade och tidskrävande karaktär. Även om den är skicklig på att underlätta smyg, är dess tillämpning i strid opraktisk, med tanke på besvärjelsens utdragna castingtid.