Det är inte ofta som en äventyrare som du blir kallad till Wizard's Keep, särskilt med så kort varsel. Du har fått brådskande nyheter från en nära vän i hållaren, som informerar dig om att de behöver personer som du själv för att skydda platsen. Det är uppenbart att någon form av leverans har ägt rum, uppenbarligen har föremålen som flyttas ett betydande värde.

Det är midsommar, men hela området är indraget i en snöstorm. Snö och is vispas upp till lakan som rullar över utsikten utanför ditt fönster, nedstigande från Deathdrop-bergen en bit bort, slingrande kring fästena i borgen som dödens kalla hand. Något stämmer inte riktigt här. Torpet ligger inom tio mil från Desert of Skulls, det borde inte finnas snö här, och absolut inte en snöstorm. Genom att låta din överaktiva fantasi vila en stund, och skylla vädret på trollkarlarna, lägger du dig i sängen och försöker ta dig till ro, faller i en störd sömn, trött från din resa till gården.

En enda ringsignal från keeps klocka signalerar början på en ny och övergiven dag... Det är midnatt. Snöplattorna fortsätter att anfalla den antika byggnaden och rikoschetterar sig från sidorna som små glassplitter. Långt borta på avstånd traskar en ensam man mot den platsen. Böjd dubbelt över sin ekkäpp spänner han ögonen i mörkret, hans lykta värdelös i detta väder. Några minuter senare når han porten.

En hög röst hörs från porthusets lyktaljus, knappt hörbar ovanför den rasande stormen.

"Sluta! I det magiska protektoratets namn, vem går dit?”

Den gamle tittar mot lyktljuset och svarar med en röst som låter ansträngd och vilsen:

"Jag är i desperat behov av skydd... kan du snälla hjälpa mig? Allt jag ber om är en säng för natten..."

Det kommer ett svar inifrån porthuset, mumlar, kvävt klagomål som frågar om besökaren är medveten om vad klockan är, när låsen klickar upp med ett högt, dovt dunk och mannen skjuts in. Flera tysta minuter senare är allt som återstår av portvakten en liten pöl av blod och pulveriserat ben som blåser runt golvet i porthuset i vinden.

Något tyst rör sig nerför korridoren som förbinder porthuset med slottets interiör. Systematiskt söker den igenom varje rum, ett efter ett. Den susar förbi dig i sömnen, till synes genom dig... och orsakar mörka och hemska mardrömmar när den passerar, och din sömn blir allt mer rastlös.
Långt senare har Something hittat sin väg till gårdens djup. Många våningar under ytan, nerför en lång korridor täckt av runor, står den framför en enorm ek- och gulddörr, bevakad av två vakter, välutbildade i magiska konster, alert och redo att avvärja attacker.
Saken susar förbi den första vakten, fortfarande inte synlig, men lämnar en känsla av rädsla och förtvivlan vart den än går.
"Deran? Är det du?"
Den första vakten tittar åt sidan och hör en röst, till synes från ingenstans, viskande och muttlande i mörkret. Innan han vet vad som händer har The Thing sugit in hans själ i magins rike. De två sekunderna av distraktion är allt som behövs för att uppnå uppgiften.
"Hej, var uppmärksam! Det är meningen att vi ska titta..."
Den andra vaktposten släpper sin vakt för en bråkdel av en sekund för att titta på den första vakten. Det han ser i vaktens plats fyller honom med fruktan och skräck. Framför honom står en sak, sammansatt av skuggor och mörker, nästan humanoid till formen, men genomskinlig som svart grumligt vatten. Tusentals omöjligt vita tänder sticker ut ur en mun som likt ebenholts, satta under två ögon, glödande röda som själva helvetets gropar, virvlande malströmmar av hat och lidande redo och hungriga att sluka. Vakten har chansen att uttala den första bråkdelen av ett enda, skräckslaget fruktansvärt skrik när hundra glittrande tentakler dyker upp ur den glupande maven, drar honom med ansiktet först in i varelsens mun och dränerar honom på hans väsen, och konsumerar på det mest smärtsamma, fruktansvärda och fruktansvärda sättet för någon dödlig varelse att avsluta sitt liv...