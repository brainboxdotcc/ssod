## Människorikets huvudstad

I hjärtat av mänskligt styre ligger den vidsträckta staden Cryptillius Centralius, placerad på en liten ö nära Great Northern Wastes längst norr om Cryptillia. Denna metropol fungerar som epicentrum där beslut ekar över hela planeten. Den mänskliga civilisationens tyglar hålls av en enastående kejsare, Haldrine IV, som utfärdar direktiv till en mängd herrar och damer som övervakar olika territorier.

Dessa herrar och damer, som uppgår till flera hundra, utövar avsevärd autonomi inom sina sfärer, eftersom kommunikationskanalerna mellan dem och kejsaren kännetecknas av plågsam långsamhet. Den förestående följden av den åldrade kejsaren Haldrine IV lägger till ett lager av komplexitet till maktdynamiken. Med kejsaren på randen att passera manteln, väntar hans många söner ivrigt på ögonblicket då en kommer att väljas till rättmätig arvinge. Denna situation förstärker inflytandet från de regionala herrarna och damerna, som för närvarande har en oöverträffad makt över mänsklighetens öde. När det politiska landskapet utvecklas, hänger Cryptillias öde i balans, format av besluten från både den centrala myndigheten och de formidabla herrarna som styr de olika länderna.

Stadens stora skala är imponerande, med höga strukturer som skrapar himlen, deras sten- och metallfasader ett bevis på mänsklighetens flitiga anda. Massiva broar sträcker sig över sammanbindande öar och skapar invecklade nätverk som underlättar flödet av människor och varor.

Arkitekturen av Cryptillius Centralius är en blandning av storhet och praktisk, med imponerande citadeller, invecklade spiror och labyrintiska befästningar som väver en komplex gobeläng mot bakgrund av det norra landskapet. Det centrala citadellet, där kejsaren bor, dominerar silhuetten, dess kolossala form är en symbol för auktoritet som är synlig från alla hörn av metropolen.

Inom stadens gränser sprider sig livliga marknader och livliga distrikt, som ekar av kadensen av olika språk och den harmoniska kulturkrocken. Gatorna är levande med ett kalejdoskop av färger, när köpmän säljer exotiska varor från avlägsna länder, och medborgare, utsmyckade i en mängd olika kläder, korsar de labyrintiska gränderna.

Cryptillius Centralius står som en ledstjärna för både styrka och bräcklighet, dess existens är beroende av den känsliga balansen mellan centraliserad auktoritet och regionala herrars autonomi. Luften bär på en påtaglig energi, laddad med spänningen av förestående succession och de ständigt närvarande ebb och flödet av politiska strömningar.

När solen går ner över Great Northern Wastes, flimrar stadens otaliga ljus till liv och förvandlar Cryptillius Centralius till en konstellation av briljans. Det är ett spektakel som fängslar fantasin, en förkroppsligande av mänsklig ambition och motståndskraft inför de vidsträckta mysterier som ligger utanför dess gränser.