## Stava: Flyga

Med hjälp av övergående flygning höjer flugbesvärjelsen kastaren till skyarna, med höjden proportionell mot deras spellcasting. Ändå finns varnande berättelser i överflöd, som berättar om fall där djärva spellcasters tappade sin flygfärdighet mitt under flygningen, och störtdyker till sin bortgång i tragiska, otidiga nedstigningar.