Orcweed, en tålig och anspråkslös växt, växer rikligt runt orcernas läger, vilket förkroppsligar motståndskraften hos den orchiska livsstilen. Trots sitt omärkliga utseende har Orcweed praktiska tillämpningar inom spellcasting. Ofta avfärdas av andra raser som enbart ogräs, Orcher inser dess värde och införlivar det i sina ritualer. När den används i trollformler, lägger Orcweed till en touch av ursprunglig styrka, och betonar den enkla och robusta karaktären hos orcisk magi. Dess förekomst nära Orc-läger gör det till en lättillgänglig resurs för dem som förstår dess underskattade potential.