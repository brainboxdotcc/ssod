## Stava: Öppna

Den öppna besvärjelsen, en huvudnyckel framkallad genom mystiska skicklighet, ger castern möjlighet att explosivt bryta upp lås och förseglade dörrar. Genom att utlösa en kontrollerad explosion i låsmekanismer och tätningar, driver denna förtrollning dörrar från deras gångjärn och klyver lådor isär. Medan det är ett mångsidigt verktyg i händerna på alla skickliga trollkastare, når dess potential sin zenit i en skicklig tjuvs kvicka fingrar. Tjuvar, skickliga i konsten att subterfight, utnyttjar Open-besvärjelsen för att reda ut hemligheter, stjäla skatter och navigera genom säkra passager med oöverträffad finess.