Desert of Skulls sträcker sig över landskapet som en ödslig och oförlåtande vidd, dess torra slätter avbryts av böljande sanddyner av fin, skiftande sand. Den obevekliga solen slår ner på den torra marken och skapar en skimrande hägring som dansar vid horisonten. Luften är tjock av den tryckande värmen, och landet verkar nästan sakna liv.

Spridda rester av forntida ruiner antyder en tid då denna öken inte var en karg ödemark. Nu reser sig dock skelettrester av sedan länge bortglömda strukturer från sanden som spöklika vaktposter, ett bevis på tidens hårda gång.

I hjärtat av denna ödslighet ligger den norra oasstaden Arrowhaven. Arrowhaven är en välkommen paus mitt i hårdheten, en bastion av liv som upprätthålls av en dold källa. Palmer vajar försiktigt i vinden, och kluster av livfull grönska ger en skarp kontrast till den omgivande öknen.

Staden är ett blygsamt men viktigt nav för resenärer som trotsar den förrädiska dödskallarnas öken. Dess arkitektur speglar både praktiska egenskaper och motståndskraft, med adobestrukturer som ger skydd mot den obevekliga solen. Smala gränder slingrar sig genom staden och erbjuder skugga och lättnad från den tryckande hettan.

Arrowhavens invånare är tåliga och fyndiga, efter att ha anpassat sig till utmaningarna med att leva i en sådan ogästvänlig miljö. Oasen fungerar som en viktig källa till vatten, och stadsborna har lärt sig att skörda dess rikedom för näring.

Trots sina tuffa omgivningar fungerar Arrowhaven som en avgörande vägpunkt för äventyrare, handlare och nomader som korsar öknen. Dess existens är ett bevis på motståndskraften hos dem som kallar det hem, och oasstaden står som en ledstjärna för liv mitt i den stora, skelettiga ödemarken i Desert of Skulls.