## Stava: Smyg

Smygbesvärjelsen, en övergående mantel av skuggor, tredubblar kastarens smygpoäng i tio stycken, vilket gör dem praktiskt taget omärkliga. Men den mystiska återstoden dröjer sig kvar, och för tre efterföljande platser efter att besvärjelsen har försvunnit, minskar kastarens smygpoäng till hälften av sitt ursprungliga värde. Skiktiga utövare av smyg måste navigera i denna dualitet försiktigt, för konsekvenserna ackumuleras med varje casting. Sådana trollformler visar sig vara oumbärliga för skurkar och infiltratörer som söker skuggorna och kringgår faran med varje steg i silhuett.