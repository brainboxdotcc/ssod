Monkgräs, ett botaniskt underverk inbäddat i de dolda hörnen av Cryptillia, har en medfödd koppling till språkens mångfaldiga gobeläng. Dess slanka, silvergröna blad svajar i harmonisk samklang med viskningarna från uråldriga tungor som bärs av osedda vindar. Örten är ofta eftersökt av både lingvister och trollkarlar, dess närvaro fungerar som en kanal för att låsa upp kommunikationens krångligheter. När det används i spellcasting, tros Monkgräs bredda sinnets mottaglighet för främmande språk, och främja en bro mellan kastaren och de språkliga mysterier som omger dem.